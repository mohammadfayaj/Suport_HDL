-- Implemnetarea metodei Quine-McCluskey
library IEEE;
use IEEE.std_logic_1164.all;

package quine_mccluskey is
end package;

package body of quine_mccluskey is
end body;
