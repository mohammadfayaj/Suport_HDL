-- Implemnetarea metodei Quine-McCluskey
library IEEE;
use IEEE.std_logic_1164.all;

package quine_mccluskey is
	
end package;

package body quine_mccluskey is
end package body;
 